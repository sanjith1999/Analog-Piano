CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 1536 451
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
24 D:\Circuit Maker\BOM.DAT
0 7
0 71 1536 451
144179218 0
0
6 Title:
5 Name:
0
0
0
24
7 Ground~
168 945 335 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 877 322 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 874 222 0 1 3
0 2
0
0 0 53360 180
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 771 338 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 433 393 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
8 Battery~
219 876 244 0 2 5
0 5 2
0
0 0 880 180
3 10V
11 -2 32 6
2 V4
15 -12 29 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
7734 0 0
0
0
8 Battery~
219 880 309 0 2 5
0 2 6
0
0 0 880 180
3 10V
11 -2 32 6
2 V3
15 -12 29 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
10 Capacitor~
219 753 313 0 2 5
0 2 8
0
0 0 848 90
5 0.61u
4 0 39 8
2 C3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
7 Ground~
168 625 207 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3549 0 0
0
0
7 Ground~
168 626 318 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 0 0 0 0
3 GND
7931 0 0
0
0
8 Battery~
219 626 298 0 2 5
0 9 10
0
0 0 880 0
4 2.4V
9 -2 37 6
2 V2
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9325 0 0
0
0
8 Battery~
219 627 238 0 2 5
0 11 2
0
0 0 880 180
4 2.4V
8 -2 36 6
2 V1
15 -12 29 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8903 0 0
0
0
10 Capacitor~
219 484 181 0 2 5
0 13 7
0
0 0 848 0
3 10n
-11 -18 10 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3834 0 0
0
0
10 Capacitor~
219 447 272 0 2 5
0 2 14
0
0 0 848 90
3 10n
11 0 32 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3363 0 0
0
0
10 Op-Amp5:A~
219 625 267 0 5 11
0 14 15 11 9 7
0
0 0 848 0
5 UA741
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 768 1 0 0 0
1 U
7668 0 0
0
0
6 AD633~
219 831 280 0 8 17
0 7 8 8 2 6 4 3 5
0
0 0 4944 0
6 AD633J
-20 -37 22 -29
2 U1
-6 -47 8 -39
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
88 0 0 256 1 0 0 0
1 U
4718 0 0
0
0
9 Resistor~
219 946 244 0 2 5
0 4 3
0
0 0 880 90
2 1k
8 0 22 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 945 292 0 3 5
0 2 4 -1
0
0 0 880 90
2 3k
8 0 22 8
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 754 273 0 2 5
0 8 7
0
0 0 880 90
2 1k
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 430 182 0 2 5
0 14 13
0
0 0 880 0
6 60.83k
-21 -14 21 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
9 Resistor~
219 385 273 0 3 5
0 2 14 -1
0
0 0 880 90
6 60.83k
-6 0 36 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 516 391 0 3 5
0 2 12 -1
0
0 0 880 0
4 100k
-14 -14 14 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 515 350 0 3 5
0 2 12 -1
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 620 361 0 2 5
0 7 12
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
31
7 2 3 0 0 4224 0 16 17 0 0 7
864 271
909 271
909 254
929 254
929 218
946 218
946 226
1 1 2 0 0 4096 0 1 18 0 0 4
945 329
945 309
945 309
945 310
6 0 4 0 0 4224 0 16 0 0 10 4
864 280
925 280
925 267
946 267
0 0 2 0 0 4096 0 0 0 5 31 2
433 369
433 328
1 0 2 0 0 8192 0 5 0 0 25 3
433 387
433 369
475 369
1 1 2 0 0 0 0 2 7 0 0 3
877 316
877 318
878 318
1 2 2 0 0 0 0 3 6 0 0 2
874 230
874 229
8 1 5 0 0 4224 0 16 6 0 0 3
864 262
874 262
874 253
5 2 6 0 0 4224 0 16 7 0 0 3
864 289
878 289
878 294
2 1 4 0 0 0 0 18 17 0 0 3
945 274
946 274
946 262
0 0 7 0 0 4096 0 0 0 26 12 3
696 218
778 218
778 255
2 1 7 0 0 0 0 19 16 0 0 3
754 255
798 255
798 262
1 0 2 0 0 0 0 4 0 0 14 2
771 332
771 332
4 1 2 0 0 8192 0 16 8 0 0 5
798 289
793 289
793 332
753 332
753 322
0 1 8 0 0 8320 0 0 19 16 0 3
787 274
787 291
754 291
3 2 8 0 0 0 0 16 16 0 0 4
798 280
787 280
787 271
798 271
2 1 8 0 0 0 0 8 19 0 0 3
753 304
754 304
754 291
1 4 9 0 0 8320 0 11 15 0 0 3
626 285
625 285
625 280
0 2 10 0 0 4224 0 0 11 0 0 2
626 318
626 309
1 3 11 0 0 4224 0 12 15 0 0 2
625 247
625 254
1 2 2 0 0 0 0 9 12 0 0 2
625 215
625 223
1 0 7 0 0 8192 0 24 0 0 26 3
638 361
681 361
681 267
2 0 12 0 0 4096 0 24 0 0 24 2
602 361
566 361
2 2 12 0 0 8320 0 22 23 0 0 4
534 391
566 391
566 350
533 350
1 1 2 0 0 0 0 23 22 0 0 4
497 350
475 350
475 391
498 391
2 5 7 0 0 4224 0 13 15 0 0 4
493 181
696 181
696 267
643 267
2 1 13 0 0 8320 0 20 13 0 0 3
448 182
448 181
475 181
0 1 14 0 0 4096 0 0 20 30 0 3
405 238
405 182
412 182
1 0 14 0 0 4224 0 15 0 0 30 4
607 261
503 261
503 238
446 238
2 2 14 0 0 0 0 21 14 0 0 4
385 255
385 238
447 238
447 263
1 1 2 0 0 8320 0 14 21 0 0 4
447 281
447 328
385 328
385 291
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2755588 1210432 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 5
0
1969190 8550464 100 100 0 0
77 66 1487 306
0 451 1536 831
211 66
208 66
1487 87
1487 186
0 0
0.0952768 0.0932624 0.204255 0.204255 1 1
12385 4
4 5 5
1
938 218
0 3 0 0 5	0 1 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
