CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
-1920 71 -384 467
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
24 D:\Circuit Maker\BOM.DAT
0 7
-1920 71 -384 467
144179219 0
0
6 Title:
5 Name:
0
0
0
20
11 Signal Gen~
195 742 174 0 64 64
0 4 2 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 -420004444
20
0 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V6
-7 -40 7 -32
0
0
29 %D %1 %2 DC 0 SIN(0 1 1k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 956 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
8 Battery~
219 956 143 0 2 5
0 6 2
0
0 0 880 0
2 12
15 -2 29 6
2 V5
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
7 Ground~
168 907 243 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
8 Battery~
219 909 190 0 2 5
0 2 7
0
0 0 880 180
2 12
12 -2 26 6
2 V4
12 -12 26 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
6 AD633~
219 855 160 0 8 17
0 5 2 4 2 7 2 3 6
0
0 0 4944 0
6 AD633J
-20 -37 22 -29
2 U2
-6 -47 8 -39
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
88 0 0 256 1 0 0 0
1 U
7734 0 0
0
0
6 Diode~
219 387 125 0 2 5
0 8 9
0
0 0 848 0
6 1N5402
-21 -18 21 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
6 DO-201
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9914 0 0
0
0
7 Ground~
168 694 295 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
7 Ground~
168 471 251 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3549 0 0
0
0
11 Signal Gen~
195 198 148 0 24 64
0 8 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1092616192 0 1073741824
0 897988541 897988541 1000593163 1036831949
20
0 10 0 2 0 1e-006 1e-006 0.005 0.1 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/2V
-15 -30 13 -22
2 V3
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 PULSE(0 2 0 1u 1u 5m 100m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
7931 0 0
0
0
7 Ground~
168 590 136 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9325 0 0
0
0
7 Ground~
168 627 254 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8903 0 0
0
0
8 Battery~
219 590 105 0 2 5
0 10 2
0
0 0 880 0
2 12
15 -2 29 6
2 V2
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3834 0 0
0
0
8 Battery~
219 629 222 0 2 5
0 2 12
0
0 0 880 180
2 12
12 -2 26 6
2 V1
12 -12 26 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3363 0 0
0
0
10 Op-Amp5:A~
219 625 170 0 5 11
0 9 11 10 12 5
0
0 0 848 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
7668 0 0
0
0
10 Capacitor~
219 443 164 0 2 5
0 2 9
0
0 0 848 90
2 1u
14 0 28 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4718 0 0
0
0
9 Resistor~
219 1064 156 0 3 5
0 2 3 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 694 270 0 3 5
0 2 11 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 694 221 0 2 5
0 11 5
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
9 Resistor~
219 518 165 0 3 5
0 2 9 -1
0
0 0 880 90
3 10k
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4871 0 0
0
0
27
1 0 2 0 0 8320 0 17 0 0 12 3
1064 174
1064 218
907 218
7 2 3 0 0 12416 0 6 17 0 0 5
888 151
923 151
923 102
1064 102
1064 138
2 0 2 0 0 0 0 1 0 0 7 2
773 179
793 179
1 3 4 0 0 12416 0 1 6 0 0 4
773 169
778 169
778 160
822 160
6 0 2 0 0 0 0 6 0 0 6 2
888 160
956 160
1 2 2 0 0 0 0 2 3 0 0 2
956 184
956 154
0 1 2 0 0 0 0 0 4 8 0 3
793 168
793 237
907 237
2 4 2 0 0 0 0 6 6 0 0 4
822 151
793 151
793 169
822 169
1 0 5 0 0 4224 0 6 0 0 19 3
822 142
694 142
694 170
1 8 6 0 0 8320 0 3 6 0 0 4
956 130
956 131
888 131
888 142
2 5 7 0 0 8320 0 5 6 0 0 3
907 175
907 169
888 169
1 1 2 0 0 0 0 4 5 0 0 2
907 237
907 199
1 1 8 0 0 4224 0 7 10 0 0 3
377 125
229 125
229 143
2 0 9 0 0 4096 0 7 0 0 25 2
397 125
443 125
1 3 10 0 0 12416 0 13 15 0 0 4
590 92
590 84
625 84
625 157
1 2 2 0 0 0 0 11 13 0 0 2
590 130
590 116
1 1 2 0 0 0 0 8 18 0 0 2
694 289
694 288
0 2 11 0 0 4224 0 0 15 20 0 4
694 245
583 245
583 176
607 176
2 5 5 0 0 128 0 19 15 0 0 3
694 203
694 170
643 170
1 2 11 0 0 0 0 19 18 0 0 2
694 239
694 252
1 0 9 0 0 0 0 15 0 0 25 4
607 164
564 164
564 122
520 122
1 0 2 0 0 0 0 9 0 0 24 2
471 245
471 222
2 0 2 0 0 128 0 10 0 0 24 4
229 153
351 153
351 222
443 222
1 1 2 0 0 0 0 16 20 0 0 4
443 173
443 222
518 222
518 183
2 2 9 0 0 8320 0 16 20 0 0 6
443 155
443 122
520 122
520 122
518 122
518 147
1 1 2 0 0 0 0 12 14 0 0 4
627 248
627 219
627 219
627 231
2 4 12 0 0 4224 0 14 15 0 0 3
627 207
627 183
625 183
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.5 0.001 0.001
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1902624 1079360 100 100 0 0
0 0 0 0
-1920 71 -1759 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 5
0
2164764 8550464 100 100 0 0
77 66 1487 696
-1920 71 -384 864
231 66
77 66
1487 127
1487 696
0 0
0.0546099 0 0.26675 -0.33 0.5 0.5
12401 0
4 0.1 5
1
1054 102
0 3 0 0 3	0 2 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
